library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CombShiftUnit is
	port();
end CombShiftUnit;